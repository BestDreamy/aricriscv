`include "define.v"

module test_reg(
    input wire[`CPU_WIDTH - 1:0] x0,
    input wire[`CPU_WIDTH - 1:0] x1,
    input wire[`CPU_WIDTH - 1:0] x2,
    input wire[`CPU_WIDTH - 1:0] x3,
    input wire[`CPU_WIDTH - 1:0] x4,
    input wire[`CPU_WIDTH - 1:0] x5,
    input wire[`CPU_WIDTH - 1:0] x6,
    input wire[`CPU_WIDTH - 1:0] x7,
    input wire[`CPU_WIDTH - 1:0] x8,
    input wire[`CPU_WIDTH - 1:0] x9,
    input wire[`CPU_WIDTH - 1:0] x10,
    input wire[`CPU_WIDTH - 1:0] x11,
    input wire[`CPU_WIDTH - 1:0] x12,
    input wire[`CPU_WIDTH - 1:0] x13,
    input wire[`CPU_WIDTH - 1:0] x14,
    input wire[`CPU_WIDTH - 1:0] x15,
    input wire[`CPU_WIDTH - 1:0] x16,
    input wire[`CPU_WIDTH - 1:0] x17,
    input wire[`CPU_WIDTH - 1:0] x18,
    input wire[`CPU_WIDTH - 1:0] x19,
    input wire[`CPU_WIDTH - 1:0] x20,
    input wire[`CPU_WIDTH - 1:0] x21,
    input wire[`CPU_WIDTH - 1:0] x22,
    input wire[`CPU_WIDTH - 1:0] x23,
    input wire[`CPU_WIDTH - 1:0] x24,
    input wire[`CPU_WIDTH - 1:0] x25,
    input wire[`CPU_WIDTH - 1:0] x26,
    input wire[`CPU_WIDTH - 1:0] x27,
    input wire[`CPU_WIDTH - 1:0] x28,
    input wire[`CPU_WIDTH - 1:0] x29,
    input wire[`CPU_WIDTH - 1:0] x30,
    input wire[`CPU_WIDTH - 1:0] x31
);
    
endmodule
